netcdf PACE_SPEXONE_OCAL.20240407T060127.L1A {
types:
  compound nomhk_dtype {
    ushort SEQCNT ;
    ushort TCPKTID ;
    ushort TCPKTSEQCTRL ;
    ubyte TCREJCODE ;
    ubyte TCFAILCODE ;
    ushort TCREJPKTID ;
    ushort TCFAILPKTID ;
    ushort TCACCCNT ;
    ushort TCREJCNT ;
    ushort TCEXECCNT ;
    ushort TCFAILCNT ;
    ushort ICUSWVER ;
    uint SYSSTATE ;
    ubyte ICUMODE ;
    ubyte EXTPPSSTAT ;
    ubyte TIMEMSGSTAT ;
    ubyte OBTSYNCSTAT ;
    ubyte MPS_ID ;
    ubyte MPS_VER ;
    ubyte EVNTCNT_DEBUG ;
    ubyte EVNTCNT_PROG ;
    ubyte EVNTCNT_WARN ;
    ubyte EVNTCNT_ERR ;
    ubyte EVNTCNT_FATAL ;
    ubyte BOOTSTATEPREV ;
    uint BOOTCNTGOOD_IM0 ;
    uint BOOTCNTGOOD_IM1 ;
    uint BOOTCNTGOOD_IM2 ;
    uint BOOTCNTGOOD_IM3 ;
    ubyte BOOTATTEMPTS_CURRIM ;
    ubyte SWIMG_LOADED ;
    ubyte SWIMG_DEFAULT ;
    ubyte SWIMG_NXTBOOT ;
    ubyte WRITEPROT ;
    ubyte BOOTCAUSE ;
    ubyte TCVER_STAT ;
    uint SPW_REG_A ;
    uint SPW_REG_B ;
    uint LAST_CRC ;
    ushort SCITM_PKTINTVL ;
    uint SCITM_BUFFREE ;
    uint64 SWEXECTIMEWC ;
    ushort ERRCNT_PLACEHOLDER_03 ;
    uint TS1_DEM_N_T ;
    uint TS2_HOUSING_N_T ;
    uint TS3_RADIATOR_N_T ;
    uint TS4_DEM_R_T ;
    uint TS5_HOUSING_R_T ;
    uint TS6_RADIATOR_R_T ;
    ushort ICU_5V_T ;
    ushort ICU_4V_T ;
    ushort ICU_HG1_T ;
    ushort ICU_HG2_T ;
    ushort ICU_MID_T ;
    ushort ICU_MCU_T ;
    ushort ICU_DIGV_T ;
    ushort ICU_4P0V_V ;
    ushort ICU_3P3V_V ;
    ushort ICU_1P2V_V ;
    ushort ICU_4P0V_I ;
    ushort ICU_3P3V_I ;
    ushort ICU_1P2V_I ;
    ubyte DEM_STATUS ;
    ubyte dummy_01 ;
    ushort ICU_5P0V_V ;
    ushort ICU_5P0V_I ;
    ubyte DEMSPWSTAT ;
    ubyte DEMRESETCNT ;
    ushort HTRGRP1_V ;
    ushort HTRGRP2_V ;
    ushort HTR1_I ;
    ushort HTR2_I ;
    ushort HTR3_I ;
    ushort HTR4_I ;
    uint HTR1_CALCPVAL ;
    uint HTR2_CALCPVAL ;
    uint HTR3_CALCPVAL ;
    uint HTR4_CALCPVAL ;
    uint HTR1_CALCIVAL ;
    uint HTR2_CALCIVAL ;
    uint HTR3_CALCIVAL ;
    uint HTR4_CALCIVAL ;
    ushort HTR1_DUTYCYCL ;
    ushort HTR2_DUTYCYCL ;
    ushort HTR3_DUTYCYCL ;
    ushort HTR4_DUTYCYCL ;
    ubyte LED1_ENADIS ;
    ubyte LED2_ENADIS ;
    uint LED1_ANODE_V ;
    uint LED1_CATH_V ;
    uint LED1_I ;
    uint LED2_ANODE_V ;
    uint LED2_CATH_V ;
    uint LED2_I ;
    uint ADC1_VCC ;
    uint ADC1_GAIN ;
    uint ADC1_REF ;
    uint ADC1_T ;
    uint ADC1_OFFSET ;
    uint ADC2_VCC ;
    uint ADC2_GAIN ;
    uint ADC2_REF ;
    uint ADC2_T ;
    uint ADC2_OFFSET ;
    ushort DEM_V ;
    ushort DEM_I ;
    ubyte REG_FW_VERSION ;
    ubyte dummy_02 ;
    ushort DET_T ;
    ubyte REG_SPW_ERROR ;
    ubyte REG_CMV_OUTOFSYNC ;
    ubyte REG_OCD_ACTUAL ;
    ubyte REG_OCD_STICKY ;
    ubyte REG_PWR_SENS ;
    ubyte REG_FLASH_STATUS ;
    ushort REG_FLASH_EDAC_BLOCK ;
  }; // nomhk_dtype
  compound science_dtype {
    ushort ICUSWVER ;
    ubyte MPS_ID ;
    ubyte MPS_VER ;
    uint TS1_DEM_N_T ;
    uint TS2_HOUSING_N_T ;
    uint TS3_RADIATOR_N_T ;
    uint TS4_DEM_R_T ;
    uint TS5_HOUSING_R_T ;
    uint TS6_RADIATOR_R_T ;
    ushort ICU_5V_T ;
    ushort ICU_4V_T ;
    ushort ICU_HG1_T ;
    ushort ICU_HG2_T ;
    ushort ICU_MID_T ;
    ushort ICU_MCU_T ;
    ushort ICU_DIGV_T ;
    ushort ICU_4P0VB_V ;
    ushort ICU_3P3V_V ;
    ushort ICU_1P2V_V ;
    ushort ICU_4P0V_I ;
    ushort ICU_3P3V_I ;
    ushort ICU_1P2V_I ;
    ushort ICU_5P0V_V ;
    ushort ICU_5P0V_I ;
    ushort DEM_V ;
    ushort DEM_I ;
    uint LED1_ANODE_V ;
    uint LED1_CATH_V ;
    uint LED1_I ;
    uint LED2_ANODE_V ;
    uint LED2_CATH_V ;
    uint LED2_I ;
    uint ADC1_VCC ;
    uint ADC1_REF ;
    uint ADC1_T ;
    uint ADC2_VCC ;
    uint ADC2_REF ;
    uint ADC2_T ;
    ubyte REG_FW_VERSION ;
    ubyte REG_NCOADDFRAMES ;
    ubyte REG_IGEN_SELECT ;
    ubyte REG_FULL_FRAME ;
    uint REG_BINNING_TABLE_START ;
    ubyte REG_CMV_OUTPUTMODE ;
    ubyte dummy_01 ;
    uint REG_COADD_BUF_START ;
    uint REG_COADD_RESA_START ;
    uint REG_COADD_RESB_START ;
    uint REG_FRAME_BUFA_START ;
    uint REG_FRAME_BUFB_START ;
    uint REG_LINE_ENABLE_START ;
    ubyte DET_REG000 ;
    ubyte dummy_02 ;
    ushort DET_NUMLINES ;
    ushort DET_START1 ;
    ushort DET_START2 ;
    ushort DET_START3 ;
    ushort DET_START4 ;
    ushort DET_START5 ;
    ushort DET_START6 ;
    ushort DET_START7 ;
    ushort DET_START8 ;
    ushort DET_NUMLINES1 ;
    ushort DET_NUMLINES2 ;
    ushort DET_NUMLINES3 ;
    ushort DET_NUMLINES4 ;
    ushort DET_NUMLINES5 ;
    ushort DET_NUMLINES6 ;
    ushort DET_NUMLINES7 ;
    ushort DET_NUMLINES8 ;
    ushort DET_SUBS ;
    ushort DET_SUBA ;
    ubyte DET_MONO ;
    ubyte DET_IMFLIP ;
    ubyte DET_EXPCNTR ;
    ubyte DET_ILVDS ;
    uint DET_EXPTIME ;
    uint DET_EXPSTEP ;
    uint DET_KP1 ;
    uint DET_KP2 ;
    ubyte DET_NOFSLOPES ;
    ubyte DET_EXPSEQ ;
    uint DET_EXPTIME2 ;
    uint DET_EXPSTEP2 ;
    ubyte DET_REG062 ;
    ubyte DET_REG063 ;
    ubyte DET_REG064 ;
    ubyte DET_REG065 ;
    ubyte DET_REG066 ;
    ubyte DET_REG067 ;
    ubyte DET_REG068 ;
    ubyte DET_EXP2_SEQ ;
    ushort DET_NOFFRAMES ;
    ubyte DET_OUTMODE ;
    ubyte DET_FOTLEN ;
    ubyte DET_ILVDSRCVR ;
    ubyte DET_REG075 ;
    ubyte DET_REG076 ;
    ubyte DET_CALIB ;
    ushort DET_TRAINPTRN ;
    uint DET_CHENA ;
    ubyte DET_ICOL ;
    ubyte DET_ICOLPR ;
    ubyte DET_IADC ;
    ubyte DET_IAMP ;
    ubyte DET_VTFL1 ;
    ubyte DET_VTFL2 ;
    ubyte DET_VTFL3 ;
    ubyte DET_VRSTL ;
    ubyte DET_REG092 ;
    ubyte DET_REG093 ;
    ubyte DET_VPRECH ;
    ubyte DET_VREF ;
    ubyte DET_REG096 ;
    ubyte DET_REG097 ;
    ubyte DET_VRAMP1 ;
    ubyte DET_VRAMP2 ;
    ushort DET_OFFSET ;
    ubyte DET_PGAGAIN ;
    ubyte DET_ADCGAIN ;
    ubyte DET_REG104 ;
    ubyte DET_REG105 ;
    ubyte DET_REG106 ;
    ubyte DET_REG107 ;
    ubyte DET_TDIG1 ;
    ubyte DET_TDIG2 ;
    ubyte DET_REG110 ;
    ubyte DET_BITMODE ;
    ubyte DET_ADCRES ;
    ubyte DET_PLLENA ;
    ubyte DET_PLLINFRE ;
    ubyte DET_PLLBYP ;
    ubyte DET_PLLRATE ;
    ubyte DET_PLLLOAD ;
    ubyte DET_DETDUM ;
    ubyte DET_REG119 ;
    ubyte DET_REG120 ;
    ubyte DET_BLACKCOL ;
    ubyte DET_REG122 ;
    ubyte DET_VBLACKSUN ;
    ubyte DET_REG124 ;
    ubyte DET_REG125 ;
    ushort DET_T ;
    ushort FTI ;
    ubyte IMDMODE ;
    ubyte dummy_03 ;
    uint IMRLEN ;
  }; // science_dtype
dimensions:
	column = 2048 ;
	hk_packets = 437 ;
	number_of_images = 1310 ;
	quaternion_elements = 4 ;
	row = 2048 ;
	samples_per_image = 203500 ;
	vector_elements = 3 ;

// global attributes:
		string :time_coverage_start = "2024-04-07T06:01:27.036" ;
		string :time_coverage_end = "2024-04-07T06:08:43.921" ;
		:processing_version = 1LL ;
		string :product_name = "PACE_SPEXONE_OCAL.20240407T060127.L1A.nc" ;
		string :date_created = "2025-08-18T11:25:08.595" ;
		string :project = "PACE Project" ;
		string :platform = "PACE" ;
		string :instrument = "SPEXone" ;
		string :title = "PACE SPEXone Level-1A Data" ;
		string :processing_level = "L1A" ;
		string :conventions = "CF-1.10, ACDD-1.3" ;
		string :standard_name_vocabulary = "CF Standard Name Table v79" ;
		string :stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		string :cdm_data_type = "swath" ;
		string :start_direction = "Ascending" ;
		string :end_direction = "Ascending" ;
		string :identifier_product_doi_authority = "https://dx.doi.org/" ;
		string :identifier_product_doi = "10.5067/PACE/SPEXONE/L1A/SCI/2" ;
		string :institution = "NASA Goddard Space Flight Center, Ocean Biology Processing Group" ;
		string :creator_name = "NASA/GSFC" ;
		string :creator_email = "data@oceancolor.gsfc.nasa.gov" ;
		string :creator_url = "https://oceancolor.gsfc.nasa.gov" ;
		string :keyword_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		string :license = "https://www.earthdata.nasa.gov/engage/open-data-services-and-software/data-and-information-policy" ;
		string :naming_authority = "gov.nasa.gsfc.sci.oceancolor" ;
		string :publisher_name = "NASA/GSFC" ;
		string :publisher_email = "data@oceancolor.gsfc.nasa.gov" ;
		string :publisher_url = "https://oceancolor.gsfc.nasa.gov" ;
		string :history = "/home/richardh/.local/bin/spx1_level01a /nfs/SPEXone/ical/archives/spx1_l0/0x12d/2024/04/07/SPX000007333.spx" ;

group: engineering_data {
  variables:
  	double HK_tlm_time(hk_packets) ;
  		string HK_tlm_time:long_name = "HK telemetry packet time" ;
  		string HK_tlm_time:description = "ICU packaging time in seconds of day" ;
  		string HK_tlm_time:calendar = "proleptic_gregorian" ;
  		HK_tlm_time:valid_min = 0. ;
  		HK_tlm_time:valid_max = 92400. ;
  		string HK_tlm_time:units = "seconds since 2024-04-07 00:00:00" ;
  	nomhk_dtype NomHK_telemetry(hk_packets) ;
  		string NomHK_telemetry:description = "An extended subset of the housekeeping parameters at 1 Hz" ;
  		string NomHK_telemetry:units = "ICU 1V2" ;
  		string NomHK_telemetry:long_name = "Sequence counter", "TC packet ID", "TC sequence control counter", "TC reject code", "TC fail code", "TC reject packet ID", "TC fail packet ID", "TC accept counter", "TC reject counter", "TC execution counter", "TC fail counter", "ICU software version", "ICU system health state", "ICU mode", "Status of external PPS", "Status time Msg", "Status of ObtSync", "MPS identifier", "MPS version", "Number of Debug events", "Number of Info/Progress events", "Number of Warning events", "Number of Error events", "Number of Fatal events", "Previous Boot State", "Amount of Im0 successful boot counts", "Amount of Im1 successful boot counts", "Amount of Im2 successful boot counts", "Amount of Im3 successful boot counts", "Number of boot attemps with current image", "Loaded and Current running SW Image", "Default SW Image", "SW Image to Load at Next Boot", "Status of Flash Write protection", "Cause of Boot", "TC verification reporting status", "Spacewire register A (host)", "Spacewire register B (DEM)", "Latest generated CRC code", "Set interval of Science TM packets (ms)", "Available free space in Science TM buffer", "Worst case SW execution time", "Error counter", "TS1 DEM nominal temperature", "TS2 housing nominal temperature", "TS3 radiator nominal temperature", "TS4 DEM redundant temperature", "TS5 housing redundant temperature", "TS6 radiator redundant temperature", "ICU 5V supply temperature", "ICU 4V supply temperature", "ICU Heater G1 supply temperature", "ICU Heater G2 supply temperature", "ICU MidBoard temperature", "ICU MCU-RAM temperature", "3v3 supply temperature", "ICU 4V bus voltage", "ICU 3.3V bus voltage", "ICU 1.2V bus voltage", "ICU 4V bus current", "ICU 3.3V bus current", "ICU 1.2V bus current", "DEM status flag", "Dummy field", "ICU 5V bus voltage", "ICU 5V bus current", "DEM spacewire status", "DEM reset counter", "Heater group 1 voltage (nominal)", "Heater group 2 voltage (redundant)", "Nominal DEM heater current", "Nominal instrument housing heater current", "Redundant DEM heater current", "Redundant instrument housing heater current", "Nominal DEM heater calculated P value", "Nominal instrument housing heater calculated P value", "Redundant DEM heater calculated P value", "Redundant instrument housing heater calculated P value", "Nominal DEM heater calculated I value", "Nominal instrument housing heater calculated I value", "Redundant DEM heater calculated I value", "Redundant instrument housing heater calculated I value", "Nominal DEM heater duty cycle", "Nominal instrument housing heater duty cycle", "Redundant DEM heater duty cycle", "Redundant instrument housing heater duty cycle", "Led 1 command enable state", "Led 2 command enable state", "Led 1 anode voltage", "Led 1 cathode voltage", "Led 1 current", "Led 2 anode voltage", "Led 2 cathode voltage", "Led 2 current", "ADC1 analog Vcc reading", "ADC1 analog gain reading", "ADC1 reference reading", "ADC1 temperature reading", "ADC1 analog offset reading", "ADC2 analog Vcc reading", "ADC2 analog gain reading", "ADC2 reference reading", "ADC2 temperature reading", "ADC2 analog offset reading", "DEM supply voltage", "DEM supply current", "DEM firmware version", "Dummy field", "Detector temperature sensor (at DEM)", "DEM spacewire error register", "Deserialize and out of sync state", "Actual OCD state", "Sticky OCD state", "Power sense enable", "EDAC error flags", "Block number with last EDAC error" ;
  	float temp_detector(hk_packets) ;
  		string temp_detector:long_name = "Detector temperature" ;
  		string temp_detector:comment = "TS1 DEM Temperature (nominal)" ;
  		string temp_detector:units = "degC" ;
  		temp_detector:valid_min = 17.83f ;
  		temp_detector:valid_max = 18.83f ;
  	float temp_housing(hk_packets) ;
  		string temp_housing:long_name = "Housekeeping temperature" ;
  		string temp_housing:comment = "TS2 Housing Temperature (nominal)" ;
  		string temp_housing:units = "degC" ;
  		temp_housing:valid_min = 19.11f ;
  		temp_housing:valid_max = 20.11f ;
  	float temp_radiator(hk_packets) ;
  		string temp_radiator:long_name = "Radiator temperature" ;
  		string temp_radiator:comment = "TS3 Radiator Temperature (nominal)" ;
  		string temp_radiator:units = "degC" ;
  		temp_radiator:valid_min = -2.f ;
  		temp_radiator:valid_max = 3.f ;
  } // group engineering_data

group: image_attributes {
  variables:
  	ubyte binning_table(number_of_images) ;
  		string binning_table:long_name = "Binning-table ID" ;
  		binning_table:valid_min = 0UB ;
  		binning_table:valid_max = 254UB ;
  	short digital_offset(number_of_images) ;
  		string digital_offset:long_name = "Digital offset" ;
  		string digital_offset:units = "1" ;
  	double exposure_time(number_of_images) ;
  		string exposure_time:long_name = "Exposure time" ;
  		string exposure_time:units = "s" ;
  	uint icu_time_sec(number_of_images) ;
  		string icu_time_sec:calendar = "tai" ;
  		icu_time_sec:valid_min = 1956528000U ;
  		icu_time_sec:valid_max = 2493072000U ;
  		string icu_time_sec:long_name = "ICU time stamp (seconds)" ;
  		string icu_time_sec:description = "Science TM parameter ICU_TIME_SEC" ;
  		string icu_time_sec:units = "seconds since 1958-01-01 00:00:00" ;
  	ushort icu_time_subsec(number_of_images) ;
  		icu_time_subsec:valid_max = 65535US ;
  		string icu_time_subsec:long_name = "ICU time stamp (sub-seconds)" ;
  		string icu_time_subsec:description = "Science TM parameter ICU_TIME_SUBSEC" ;
  		string icu_time_subsec:units = "1/65536 seconds" ;
  		icu_time_subsec:valid_min = 0US ;
  	uint image_id(number_of_images) ;
  		string image_id:long_name = "Image counter from power-up" ;
  		image_id:valid_min = 0U ;
  		image_id:valid_max = 16383U ;
  	double image_time(number_of_images) ;
  		string image_time:long_name = "Image time" ;
  		string image_time:description = "Integration start time in seconds of day" ;
  		string image_time:calendar = "proleptic_gregorian" ;
  		image_time:valid_min = 0. ;
  		image_time:valid_max = 92400. ;
  		string image_time:units = "seconds since 2024-04-07 00:00:00" ;
  	ushort nr_coadditions(number_of_images) ;
  		string nr_coadditions:units = "1" ;
  		string nr_coadditions:long_name = "Number of coadditions" ;
  		nr_coadditions:valid_min = 1US ;
  	double timedelta_centre(number_of_images) ;
  		string timedelta_centre:description = "Add this offset to image-time (MPS specific)" ;
  		string timedelta_centre:units = "s" ;
  		string timedelta_centre:long_name = "Time-delta to centre of integration time" ;
  } // group image_attributes

group: navigation_data {
  dimensions:
  	att_time = UNLIMITED ; // (0 currently)
  	orb_time = UNLIMITED ; // (0 currently)
  	tilt_time = UNLIMITED ; // (0 currently)
  variables:
  	float att_quat(att_time, quaternion_elements) ;
  		string att_quat:long_name = "Attitude quaternions (J2000 to spacecraft)" ;
  		string att_quat:units = "seconds" ;
  		att_quat:valid_min = -1.f ;
  		att_quat:valid_max = 1.f ;
  	float att_rate(att_time, vector_elements) ;
  		string att_rate:long_name = "Attitude angular rates in spacecraft frame" ;
  		string att_rate:units = "radians/second" ;
  		att_rate:valid_min = -0.004f ;
  		att_rate:valid_max = 0.004f ;
  	double att_time(att_time) ;
  		string att_time:long_name = "Attitude sample time (seconds of day)" ;
  		string att_time:units = "seconds since %Y-%m-%d %H:%M:%S" ;
  		string att_time:calendar = "proleptic_gregorian" ;
  		att_time:valid_min = 0. ;
  		att_time:valid_max = 92400. ;
  	uint64 coverage_quality ;
  		string coverage_quality:long_name = "Coverage quality of attitude data" ;
  		string coverage_quality:standard_name = "status_flag" ;
  		coverage_quality:valid_range = 0LL, 15LL ;
  		coverage_quality:flag_values = 0LL, 1LL, 2LL, 4LL, 8LL ;
  		string coverage_quality:flag_meanings = "good missing-samples too_short_extends no_extend_at_start no_extend_at_end" ;
  	float orb_alt(orb_time) ;
  		orb_alt:valid_max = 710000.f ;
  		string orb_alt:long_name = "Orbit altitude" ;
  		string orb_alt:units = "meters" ;
  		orb_alt:valid_min = 670000.f ;
  	float orb_lat(orb_time) ;
  		string orb_lat:units = "degrees_north" ;
  		orb_lat:valid_min = -90.f ;
  		string orb_lat:long_name = "Orbit latitude (degrees North)" ;
  		orb_lat:valid_max = 90.f ;
  	float orb_lon(orb_time) ;
  		orb_lon:valid_max = 180.f ;
  		string orb_lon:long_name = "Orbit longitude (degrees East)" ;
  		string orb_lon:units = "degrees_east" ;
  		orb_lon:valid_min = -180.f ;
  	float orb_pos(orb_time, vector_elements) ;
  		string orb_pos:long_name = "Orbit position vectors (ECR)" ;
  		string orb_pos:units = "meters" ;
  		orb_pos:valid_min = -7200000.f ;
  		orb_pos:valid_max = 7200000.f ;
  	double orb_time(orb_time) ;
  		string orb_time:long_name = "Orbit vector time (seconds of day)" ;
  		string orb_time:calendar = "proleptic_gregorian" ;
  		string orb_time:units = "seconds since %Y-%m-%d %H:%M:%S" ;
  		orb_time:valid_min = 0. ;
  		orb_time:valid_max = 92400. ;
  	float orb_vel(orb_time, vector_elements) ;
  		string orb_vel:long_name = "Orbit velocity vectors (ECR)" ;
  		string orb_vel:units = "meters/second" ;
  		orb_vel:valid_min = -7600.f ;
  		orb_vel:valid_max = 7600.f ;
  	float tilt(tilt_time) ;
  		string tilt:long_name = "Tilt angle" ;
  		string tilt:units = "degrees" ;
  		tilt:valid_min = -20.1f ;
  		tilt:valid_max = 20.1f ;
  	ubyte tilt_flag(tilt_time) ;
  		string tilt_flag:flag_meanings = "Valid Not_initialized" ;
  		string tilt_flag:long_name = "Tilt quality flag" ;
  		tilt_flag:flag_values = 0UB, 1UB ;
  	double tilt_time(tilt_time) ;
  		string tilt_time:long_name = "Tilt sample time (seconds of day)" ;
  		string tilt_time:calendar = "proleptic_gregorian" ;
  		string tilt_time:units = "seconds since %Y-%m-%d %H:%M:%S" ;
  		tilt_time:valid_min = 0. ;
  		tilt_time:valid_max = 92400. ;
  } // group navigation_data

group: processing_control {

  // group attributes:
  		string :software_name = "spx1_level01a" ;
  		string :software_version = "1.4.18.dev24" ;
  		string :software_description = "SPEXone L0-L1A processor (SRON)" ;
  		string :software_url = "https://github.com/rmvanhees/pyspex" ;
  		string :software_doi = "https://doi.org/10.5281/zenodo.5705691" ;

  group: input_parameters {

    // group attributes:
    		string :outdir = "/data/richardh/git/pyspex" ;
    		string :outfile = "" ;
    		string :debug = "False" ;
    		string :dump = "False" ;
    		string :verbose = "30" ;
    		string :compression = "False" ;
    		string :processing_version = "1" ;
    		string :eclipse = "None" ;
    		string :yaml_fl = "None" ;
    		string :hkt_list = "" ;
    		string :l0_format = "dsb" ;
    		string :l0_list = "SPX000007333.spx" ;
    } // group input_parameters
  } // group processing_control

group: science_data {
  variables:
  	ushort detector_images(number_of_images, samples_per_image) ;
  		string detector_images:long_name = "Detector pixel values" ;
  		string detector_images:units = "counts" ;
  		detector_images:valid_min = 0US ;
  		detector_images:valid_max = 65534US ;
  	science_dtype science_hk(number_of_images) ;
  		string science_hk:comment = "a subset of DemHK and NomHK parameters" ;
  		string science_hk:units = "ICU 1V2", "DEM internal generator register (0=test generator", "DEM frame mode register (1=diagnostic", "Number of active LVDS channels (1=science (8 ch)", "Digital offset", "Frame Trigger Interval", "Image data mode (0=DEM" ;
  		string science_hk:long_name = "ICU software version", "MPS identifier", "MPS version", "TS1 DEM nominal temperature", "TS2 housing nominal temperature", "TS3 radiator nominal temperature", "TS4 DEM redundant temperature", "TS5 housing redundant temperature", "TS6 radiator redundant temperature", "ICU 5V supply temperature", "ICU 4V supply temperature", "ICU Heater G1 supply temperature", "ICU Heater G2 supply temperature", "ICU MidBoard temperature", "ICU MCU-RAM temperature", "3v3 supply temperature", "ICU 4V bus voltage", "ICU 3.3V bus voltage", "ICU 1.2V bus voltage", "ICU 4V bus current", "ICU 3.3V bus current", "ICU 1.2V bus current", "ICU 5V bus voltage", "ICU 5V bus current", "DEM supply voltage", "DEM supply current", "Led 1 measured anode voltage", "Led 1 measured cathode voltage", "Led 1 measured current", "Led 2 measured anode voltage", "Led 2 measured cathode voltage", "Led 2 measured current", "ADC1 analog Vcc reading", "ADC1 reference reading", "ADC1 temperature reading", "ADC2 analog Vcc reading", "ADC2 reference reading", "ADC2 temperature reading", "DEM firmware version register", "DEM co-adding register", "1=detector)", "2=science)", "Start address of applicable binning table", "3=diagnostic (2 ch))", "Dummy field", "Address of co-adder buffer (intermediate)", "Address of coadding buffer A (final)", "Address of coadding buffer B (final)", "Address of buffer A (binned)", "Address of buffer B (binned)", "Address of line-enabling table", "Detector register 000 content", "Dummy field", "Number of rows read-out by sensor", "Offset in rows (block 1)", "Offset in rows (block 2)", "Offset in rows (block 3)", "Offset in rows (block 4)", "Offset in rows (block 5)", "Offset in rows (block 6)", "Offset in rows (block 7)", "Offset in rows (block 8)", "Number of rows read-out by sensor (block 1)", "Number of rows read-out by sensor (block 2)", "Number of rows read-out by sensor (block 3)", "Number of rows read-out by sensor (block 4)", "Number of rows read-out by sensor (block 5)", "Number of rows read-out by sensor (block 6)", "Number of rows read-out by sensor (block 7)", "Number of rows read-out by sensor (block 8)", "Number of rows to skip", "Number of rows to skip", "Monochrome sensor", "Image flipping", "Bits for INTE_SYNC", "LVDS current", "Exposure time", "Step size for increasing exposure times", "t$_{exp}$ at kneepoint 1 (not used)", "t$_{exp}$ at kneepoint 2 (not used)", "Number of slopes (piecewise linear response)", "Number of frames in multi-frame mode", "Exposure time (seconds)", "Step size for increasing exposure times", "Detector register 062 content", "Detector register 063 content", "Detector register 064 content", "Detector register 065 content", "Detector register 066 content", "Detector register 067 content", "Detector register 068 content", "Number of frames in multi-frame mode", "Number of frames grabbed and sent by sensor", "Number of LVDS interfaces (1=8 ch or 3=2 ch)", "Frame overhead time", "Current LVDS receiver", "Detector register 075 content", "Detector register 076 content", "Parameters COL_calib and ADC_calib", "Training pattern", "Enable/Disable channels to save power", "I$_{col}$", "I$_{col_prech}$", "I$_{ADC}$", "I$_{amp}$", "V$_{low1}$", "V$_{low2}$", "V$_{low3}$", "V$_{res_low}$", "Detector register 092 content", "Detector register 093 content", "V$_{prech}$", "V$_{ref}$", "Detector register 000 content", "Detector register 000 content", "Voltage first ramp", "Voltage second ramp", "dark-level = 70 + Offset", "Analog gain by PGA (first bit BLACKCOL)", "Digital gain by ADC", "Detector register 104 content", "Detector register 105 content", "Detector register 106 content", "Detector register 107 content", "Detector register 108 content", "Detector register 109 content", "Detector register 110 content", "Bits per pixel (default 10)", "Bits per pixel (default 10)", "Status internal PLL", "PLL input frequency", "Use or bypass internal PLL", "Set to 9 in case of 10 bit mode", "Set to 8 in case of 10 bit mode", "Dummy", "Detector register 119 content", "Detector register 120 content", "Put first 16 columns to a black reference", "Detector register 122 content", "V$_{blacksun}$", "Detector register 124 content", "Detector register 125 content", "Detector temperature sensor (at DEM)", "LSB=0.1 ms (science=667 or 15 Hz)", "1=ICU test generator)", "Dummy field", "Size of image data in bytes" ;
  } // group science_data
}
