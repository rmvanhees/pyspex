netcdf PACE_SPEXONE.20240701T055831.L1A {
types:
  compound science_dtype {
    ushort ICUSWVER ;
    ubyte MPS_ID ;
    ubyte MPS_VER ;
    uint TS1_DEM_N_T ;
    uint TS2_HOUSING_N_T ;
    uint TS3_RADIATOR_N_T ;
    uint TS4_DEM_R_T ;
    uint TS5_HOUSING_R_T ;
    uint TS6_RADIATOR_R_T ;
    short ICU_5V_T ;
    short ICU_4V_T ;
    short ICU_HG1_T ;
    short ICU_HG2_T ;
    short ICU_MID_T ;
    short ICU_MCU_T ;
    short ICU_DIGV_T ;
    ushort ICU_4P0V_V ;
    ushort ICU_3P3V_V ;
    ushort ICU_1P2V_V ;
    ushort ICU_4P0V_I ;
    ushort ICU_3P3V_I ;
    ushort ICU_1P2V_I ;
    ushort ICU_5P0V_V ;
    ushort ICU_5P0V_I ;
    ushort DEM_V ;
    ushort DEM_I ;
    uint LED1_ANODE_V ;
    uint LED1_CATH_V ;
    uint LED1_I ;
    uint LED2_ANODE_V ;
    uint LED2_CATH_V ;
    uint LED2_I ;
    uint ADC1_VCC ;
    uint ADC1_REF ;
    uint ADC1_T ;
    uint ADC2_VCC ;
    uint ADC2_REF ;
    uint ADC2_T ;
    ubyte REG_FW_VERSION ;
    ubyte REG_NCOADDFRAMES ;
    ubyte REG_IGEN_SELECT ;
    ubyte REG_FULL_FRAME ;
    uint REG_BINNING_TABLE_START ;
    ubyte REG_CMV_OUTPUTMODE ;
    ubyte dummy_01 ;
    uint REG_COADD_BUF_START ;
    uint REG_COADD_RESA_START ;
    uint REG_COADD_RESB_START ;
    uint REG_FRAME_BUFA_START ;
    uint REG_FRAME_BUFB_START ;
    uint REG_LINE_ENABLE_START ;
    ubyte DET_REG000 ;
    ubyte dummy_02 ;
    ushort DET_NUMLINES ;
    ushort DET_START1 ;
    ushort DET_START2 ;
    ushort DET_START3 ;
    ushort DET_START4 ;
    ushort DET_START5 ;
    ushort DET_START6 ;
    ushort DET_START7 ;
    ushort DET_START8 ;
    ushort DET_NUMLINES1 ;
    ushort DET_NUMLINES2 ;
    ushort DET_NUMLINES3 ;
    ushort DET_NUMLINES4 ;
    ushort DET_NUMLINES5 ;
    ushort DET_NUMLINES6 ;
    ushort DET_NUMLINES7 ;
    ushort DET_NUMLINES8 ;
    ushort DET_SUBS ;
    ushort DET_SUBA ;
    ubyte DET_MONO ;
    ubyte DET_IMFLIP ;
    ubyte DET_EXPCNTR ;
    ubyte DET_ILVDS ;
    uint DET_EXPTIME ;
    uint DET_EXPSTEP ;
    uint DET_KP1 ;
    uint DET_KP2 ;
    ubyte DET_NOFSLOPES ;
    ubyte DET_EXPSEQ ;
    uint DET_EXPTIME2 ;
    uint DET_EXPSTEP2 ;
    ubyte DET_REG062 ;
    ubyte DET_REG063 ;
    ubyte DET_REG064 ;
    ubyte DET_REG065 ;
    ubyte DET_REG066 ;
    ubyte DET_REG067 ;
    ubyte DET_REG068 ;
    ubyte DET_EXP2_SEQ ;
    ushort DET_NOFFRAMES ;
    ubyte DET_OUTMODE ;
    ubyte DET_FOTLEN ;
    ubyte DET_ILVDSRCVR ;
    ubyte DET_REG075 ;
    ubyte DET_REG076 ;
    ubyte DET_CALIB ;
    ushort DET_TRAINPTRN ;
    uint DET_CHENA ;
    ubyte DET_ICOL ;
    ubyte DET_ICOLPR ;
    ubyte DET_IADC ;
    ubyte DET_IAMP ;
    ubyte DET_VTFL1 ;
    ubyte DET_VTFL2 ;
    ubyte DET_VTFL3 ;
    ubyte DET_VRSTL ;
    ubyte DET_REG092 ;
    ubyte DET_REG093 ;
    ubyte DET_VPRECH ;
    ubyte DET_VREF ;
    ubyte DET_REG096 ;
    ubyte DET_REG097 ;
    ubyte DET_VRAMP1 ;
    ubyte DET_VRAMP2 ;
    ushort DET_OFFSET ;
    ubyte DET_PGAGAIN ;
    ubyte DET_ADCGAIN ;
    ubyte DET_REG104 ;
    ubyte DET_REG105 ;
    ubyte DET_REG106 ;
    ubyte DET_REG107 ;
    ubyte DET_TDIG1 ;
    ubyte DET_TDIG2 ;
    ubyte DET_REG110 ;
    ubyte DET_BITMODE ;
    ubyte DET_ADCRES ;
    ubyte DET_PLLENA ;
    ubyte DET_PLLINFRE ;
    ubyte DET_PLLBYP ;
    ubyte DET_PLLRATE ;
    ubyte DET_PLLLOAD ;
    ubyte DET_DETDUM ;
    ubyte DET_REG119 ;
    ubyte DET_REG120 ;
    ubyte DET_BLACKCOL ;
    ubyte DET_REG122 ;
    ubyte DET_VBLACKSUN ;
    ubyte DET_REG124 ;
    ubyte DET_REG125 ;
    ushort DET_T ;
    ushort FTI ;
    ubyte IMDMODE ;
    ubyte dummy_03 ;
    uint IMRLEN ;
  }; // science_dtype
  compound nomhk_dtype {
    ushort SEQCNT ;
    ushort TCPKTID ;
    ushort TCPKTSEQCTRL ;
    ubyte TCREJCODE ;
    ubyte TCFAILCODE ;
    ushort TCREJPKTID ;
    ushort TCFAILPKTID ;
    ushort TCACCCNT ;
    ushort TCREJCNT ;
    ushort TCEXECCNT ;
    ushort TCFAILCNT ;
    ushort ICUSWVER ;
    uint SYSSTATE ;
    ubyte ICUMODE ;
    ubyte EXTPPSSTAT ;
    ubyte TIMEMSGSTAT ;
    ubyte OBTSYNCSTAT ;
    ubyte MPS_ID ;
    ubyte MPS_VER ;
    ubyte EVNTCNT_DEBUG ;
    ubyte EVNTCNT_PROG ;
    ubyte EVNTCNT_WARN ;
    ubyte EVNTCNT_ERR ;
    ubyte EVNTCNT_FATAL ;
    ubyte BOOTSTATEPREV ;
    uint BOOTCNTGOOD_IM0 ;
    uint BOOTCNTGOOD_IM1 ;
    uint BOOTCNTGOOD_IM2 ;
    uint BOOTCNTGOOD_IM3 ;
    ubyte BOOTATTEMPTS_CURRIM ;
    ubyte MPS_ACT_STATUS ;
    ubyte SWIMG_LOADED ;
    ubyte SWIMG_DEFAULT ;
    ubyte SWIMG_NXTBOOT ;
    ubyte WRITEPROT ;
    ubyte BOOTCAUSE ;
    ubyte TCVER_STAT ;
    uint SPW_REG_A ;
    uint SPW_REG_B ;
    uint LAST_CRC ;
    ushort SCITM_PKTINTVL ;
    uint SCITM_BUFFREE ;
    uint64 SWEXECTIMEWC ;
    ushort ERRCNT_PLACEHOLDER_03 ;
    uint TS1_DEM_N_T ;
    uint TS2_HOUSING_N_T ;
    uint TS3_RADIATOR_N_T ;
    uint TS4_DEM_R_T ;
    uint TS5_HOUSING_R_T ;
    uint TS6_RADIATOR_R_T ;
    ushort ICU_5V_T ;
    ushort ICU_4V_T ;
    ushort ICU_HG1_T ;
    ushort ICU_HG2_T ;
    ushort ICU_MID_T ;
    ushort ICU_MCU_T ;
    ushort ICU_DIGV_T ;
    ushort ICU_4P0V_V ;
    ushort ICU_3P3V_V ;
    ushort ICU_1P2V_V ;
    ushort ICU_4P0V_I ;
    ushort ICU_3P3V_I ;
    ushort ICU_1P2V_I ;
    ubyte DEM_STATUS ;
    ubyte dummy_01 ;
    ushort ICU_5P0V_V ;
    ushort ICU_5P0V_I ;
    ubyte DEMSPWSTAT ;
    ubyte DEMRESETCNT ;
    ushort HTRGRP1_V ;
    ushort HTRGRP2_V ;
    ushort HTR1_I ;
    ushort HTR2_I ;
    ushort HTR3_I ;
    ushort HTR4_I ;
    float HTR1_CALCPVAL ;
    float HTR2_CALCPVAL ;
    float HTR3_CALCPVAL ;
    float HTR4_CALCPVAL ;
    float HTR1_CALCIVAL ;
    float HTR2_CALCIVAL ;
    float HTR3_CALCIVAL ;
    float HTR4_CALCIVAL ;
    ushort HTR1_DUTYCYCL ;
    ushort HTR2_DUTYCYCL ;
    ushort HTR3_DUTYCYCL ;
    ushort HTR4_DUTYCYCL ;
    ubyte LED1_ENADIS ;
    ubyte LED2_ENADIS ;
    uint LED1_ANODE_V ;
    uint LED1_CATH_V ;
    uint LED1_I ;
    uint LED2_ANODE_V ;
    uint LED2_CATH_V ;
    uint LED2_I ;
    uint ADC1_VCC ;
    uint ADC1_GAIN ;
    uint ADC1_REF ;
    uint ADC1_T ;
    uint ADC1_OFFSET ;
    uint ADC2_VCC ;
    uint ADC2_GAIN ;
    uint ADC2_REF ;
    uint ADC2_T ;
    uint ADC2_OFFSET ;
    ushort DEM_V ;
    ushort DEM_I ;
    ubyte REG_FW_VERSION ;
    ubyte dummy_02 ;
    ushort DET_T ;
    ubyte REG_SPW_ERROR ;
    ubyte REG_CMV_OUTOFSYNC ;
    ubyte REG_OCD_ACTUAL ;
    ubyte REG_OCD_STICKY ;
    ubyte REG_PWR_SENS ;
    ubyte REG_FLASH_STATUS ;
    ushort REG_FLASH_EDAC_BLOCK ;
    uint SW_MAIN_LOOP_COUNT ;
  }; // nomhk_dtype
dimensions:
	number_of_images = 8669 ;
	samples_per_image = 203500 ;
	hk_packets = 2907 ;
variables:
	string processor_configuration ;
		processor_configuration:comment = "Configuration parameters used during the processor run that produced this file." ;
		processor_configuration:markup_language = "YAML" ;

// global attributes:
		:creator_name = "NASA/GSFC" ;
		:creator_email = "data@oceancolor.gsfc.nasa.gov" ;
		:creator_url = "http://oceancolor.gsfc.nasa.gov" ;
		:institution = "NASA Goddard Space Flight Center, Ocean Biology Processing Group" ;
		:publisher_name = "NASA/GSFC" ;
		:publisher_email = "data@oceancolor.gsfc.nasa.gov" ;
		:publisher_url = "http://oceancolor.gsfc.nasa.gov" ;
		:standard_name_vocabulary = "CF Standard Name Table v79" ;
		:keyword_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:license = "http://science.nasa.gov/earth-science/earth-science-data/data-information-policy/" ;
		:naming_authority = "gov.nasa.gsfc.sci.oceancolor" ;
		:project = "PACE Project" ;
		:conventions = "CF-1.8 ACDD-1.3" ;
		:title = "PACE SPEXone Level-1A Data" ;
		:instrument = "SPEXone" ;
		:platform = "PACE" ;
		:stdname_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:processing_level = "L1A" ;
		:cdm_data_type = "swath" ;
		:product_name = "PACE_SPEXONE.20240701T055831.L1A.nc" ;
		:start_direction = "Ascending" ;
		:end_direction = "Ascending" ;
		:time_coverage_start = "2024-07-01T05:58:31.606" ;
		:time_coverage_end = "2024-07-01T06:46:53.319" ;
		:processing_version = 1LL ;
		:identifier_product_doi_authority = "http://dx.doi.org/" ;
		:identifier_product_doi = "10.5067/PACE/SPEXONE/L1A/SCI/2" ;
		:date_created = "2024-08-14T11:45:37.748" ;
		:history = "/home/richardh/.local/bin/spx1_level01a --verbose info --yaml examples/l1agen_spex/run_20240701055800.yaml" ;

group: image_attributes {
  variables:
  	uint icu_time_sec(number_of_images) ;
  		icu_time_sec:long_name = "ICU time stamp (seconds)" ;
  		icu_time_sec:description = "Science TM parameter ICU_TIME_SEC." ;
  		icu_time_sec:valid_min = 1956528000U ;
  		icu_time_sec:valid_max = 2493072000U ;
  		icu_time_sec:units = "seconds since 1958-01-01 00:00:00 TAI" ;
  	ushort icu_time_subsec(number_of_images) ;
  		icu_time_subsec:long_name = "ICU time stamp (sub-seconds)" ;
  		icu_time_subsec:description = "Science TM parameter ICU_TIME_SUBSEC." ;
  		icu_time_subsec:valid_min = 0US ;
  		icu_time_subsec:valid_max = 65535US ;
  		icu_time_subsec:units = "1/65536 s" ;
  	double image_time(number_of_images) ;
  		image_time:_FillValue = -32767. ;
  		image_time:long_name = "image time" ;
  		image_time:description = "Integration start time in seconds of day." ;
  		image_time:units = "seconds since 2024-07-01 00:00:00" ;
  		image_time:year = "2024" ;
  		image_time:month = "7" ;
  		image_time:day = "1" ;
  		image_time:valid_min = 0. ;
  		image_time:valid_max = 92304. ;
  	double timedelta_centre(number_of_images) ;
  		timedelta_centre:_FillValue = -32767. ;
  		timedelta_centre:long_name = "time-delta to centre of integration time" ;
  		timedelta_centre:description = "Add this offset to image-time (MPS specific)." ;
  		timedelta_centre:units = "s" ;
  	ushort nr_coadditions(number_of_images) ;
  		nr_coadditions:_FillValue = 0US ;
  		nr_coadditions:long_name = "number of coadditions" ;
  		nr_coadditions:valid_min = 1US ;
  		nr_coadditions:units = "1" ;
  	double exposure_time(number_of_images) ;
  		exposure_time:_FillValue = 0. ;
  		exposure_time:long_name = "exposure time" ;
  		exposure_time:units = "s" ;
  	int image_ID(number_of_images) ;
  		image_ID:long_name = "image counter from power-up" ;
  		image_ID:valid_min = 0 ;
  		image_ID:valid_max = 2147483647 ;
  	ubyte binning_table(number_of_images) ;
  		binning_table:long_name = "binning-table ID" ;
  		binning_table:valid_min = 0UB ;
  		binning_table:valid_max = 255UB ;
  	short digital_offset(number_of_images) ;
  		digital_offset:long_name = "digital offset" ;
  		digital_offset:units = "1" ;
  } // group image_attributes

group: science_data {
  variables:
  	ushort detector_images(number_of_images, samples_per_image) ;
  		detector_images:_FillValue = 65535US ;
  		detector_images:long_name = "detector pixel values" ;
  		detector_images:valid_min = 0US ;
  		detector_images:valid_max = 65534US ;
  		detector_images:units = "counts" ;
  	science_dtype detector_telemetry(number_of_images) ;
  		detector_telemetry:long_name = "SPEX science telemetry" ;
  		detector_telemetry:comment = "A subset of MPS and housekeeping parameters." ;
  } // group science_data

group: engineering_data {
  variables:
  	double HK_tlm_time(hk_packets) ;
  		HK_tlm_time:_FillValue = -32767. ;
  		HK_tlm_time:long_name = "HK telemetry packet time" ;
  		HK_tlm_time:description = "Packaging time in seconds of day." ;
  		HK_tlm_time:units = "seconds since 2024-07-01 00:00:00" ;
  		HK_tlm_time:year = "2024" ;
  		HK_tlm_time:month = "7" ;
  		HK_tlm_time:day = "1" ;
  		HK_tlm_time:valid_min = 0. ;
  		HK_tlm_time:valid_max = 92304. ;
  	nomhk_dtype NomHK_telemetry(hk_packets) ;
  		NomHK_telemetry:long_name = "SPEX nominal-HK telemetry" ;
  		NomHK_telemetry:comment = "An extended subset of the housekeeping parameters." ;
  	float temp_detector(hk_packets) ;
  		temp_detector:long_name = "detector temperature" ;
  		temp_detector:comment = "TS1 DEM Temperature (nominal)." ;
  		temp_detector:valid_min = 17.83f ;
  		temp_detector:valid_max = 18.83f ;
  		temp_detector:units = "degC" ;
  	float temp_housing(hk_packets) ;
  		temp_housing:long_name = "housing temperature" ;
  		temp_housing:comment = "TS2 Housing Temperature (nominal)." ;
  		temp_housing:valid_min = 19.11f ;
  		temp_housing:valid_max = 20.11f ;
  		temp_housing:units = "degC" ;
  	float temp_radiator(hk_packets) ;
  		temp_radiator:long_name = "radiator temperature" ;
  		temp_radiator:comment = "TS3 Radiator Temperature (nominal)." ;
  		temp_radiator:valid_min = -2.f ;
  		temp_radiator:valid_max = 3.f ;
  		temp_radiator:units = "degC" ;
  } // group engineering_data

group: processing_control {

  // group attributes:
  		:software_name = "spx1_level01a" ;
  		:software_description = "SPEXone L0-L1A processor (SRON)" ;
  		:software_url = "https://github.com/rmvanhees/pyspex" ;
  		:software_version = "1.4.14.dev15" ;
  		:software_doi = "https://doi.org/10.5281/zenodo.5705691" ;
  		:icu_sw_version = "0x12d" ;

  group: input_parameters {

    // group attributes:
    		:debug = "False" ;
    		:dump = "False" ;
    		:verbose = "20" ;
    		:compression = "False" ;
    		:outdir = "L1A" ;
    		:outfile = "" ;
    		:processing_version = "1" ;
    		:eclipse = "False" ;
    		:yaml_fl = "examples/l1agen_spex/run_20240701055800.yaml" ;
    		:hkt_list = "PACE.20240701T055223.HKT.nc,PACE.20240701T055757.HKT.nc,PACE.20240701T060332.HKT.nc,PACE.20240701T060908.HKT.nc,PACE.20240701T061445.HKT.nc,PACE.20240701T062022.HKT.nc,PACE.20240701T062600.HKT.nc,PACE.20240701T063137.HKT.nc,PACE.20240701T063714.HKT.nc,PACE.20240701T064252.HKT.nc" ;
    		:l0_format = "dsb" ;
    		:l0_list = "SPX000016243.spx,SPX000016244.spx,SPX000016245.spx,SPX000016246.spx,SPX000016247.spx,SPX000016248.spx,SPX000016249.spx" ;
    } // group input_parameters
  } // group processing_control

group: navigation_data {
  dimensions:
  	att_time = 2921 ;
  	quaternion_elements = 4 ;
  	vector_elements = 3 ;
  	orb_time = 730 ;
  	tilt_time = 2923 ;
  variables:
  	double att_time(att_time) ;
  		att_time:long_name = "Attitude sample time (seconds of day)" ;
  		att_time:valid_max = 172800. ;
  		att_time:calendar = "proleptic_gregorian" ;
  		att_time:_FillValue = -32767. ;
  		att_time:units = "seconds since 2024-07-01" ;
  		att_time:valid_min = 0. ;
  	float att_quat(att_time, quaternion_elements) ;
  		att_quat:units = "seconds" ;
  		att_quat:_FillValue = -32767.f ;
  		att_quat:long_name = "Attitude quaternions (J2000 to spacecraft)" ;
  		att_quat:valid_min = -1.f ;
  		att_quat:valid_max = 1.f ;
  	float att_rate(att_time, vector_elements) ;
  		att_rate:_FillValue = -32767.f ;
  		att_rate:long_name = "Attitude angular rates in spacecraft frame" ;
  		att_rate:valid_min = -0.004f ;
  		att_rate:valid_max = 0.004f ;
  		att_rate:units = "radians/second" ;
  	double orb_time(orb_time) ;
  		orb_time:long_name = "Orbit vector time (seconds of day)" ;
  		orb_time:valid_max = 172800. ;
  		orb_time:calendar = "proleptic_gregorian" ;
  		orb_time:_FillValue = -32767. ;
  		orb_time:units = "seconds since 2024-07-01" ;
  		orb_time:valid_min = 0. ;
  	float orb_pos(orb_time, vector_elements) ;
  		orb_pos:units = "meters" ;
  		orb_pos:_FillValue = -9999999.f ;
  		orb_pos:long_name = "Orbit position vectors (ECR)" ;
  		orb_pos:valid_min = -7200000.f ;
  		orb_pos:valid_max = 7200000.f ;
  	float orb_vel(orb_time, vector_elements) ;
  		orb_vel:_FillValue = -32767.f ;
  		orb_vel:long_name = "Orbit velocity vectors (ECR)" ;
  		orb_vel:valid_min = -7600.f ;
  		orb_vel:valid_max = 7600.f ;
  		orb_vel:units = "meters/second" ;
  	double orb_lon(orb_time) ;
  		orb_lon:_FillValue = -32767. ;
  		orb_lon:long_name = "Orbit longitude (degrees East)" ;
  		orb_lon:valid_min = -180. ;
  		orb_lon:valid_max = 180. ;
  		orb_lon:units = "degrees_east" ;
  	double orb_lat(orb_time) ;
  		orb_lat:_FillValue = -32767. ;
  		orb_lat:long_name = "Orbit latitude (degrees North)" ;
  		orb_lat:valid_min = -90. ;
  		orb_lat:valid_max = 90. ;
  		orb_lat:units = "degrees_north" ;
  	double orb_alt(orb_time) ;
  		orb_alt:_FillValue = -32767. ;
  		orb_alt:long_name = "Orbit altitude" ;
  		orb_alt:units = "meters" ;
  		orb_alt:valid_min = 670000. ;
  		orb_alt:valid_max = 710000. ;
  	double tilt_time(tilt_time) ;
  		tilt_time:long_name = "Tilt sample time (seconds of day)" ;
  		tilt_time:valid_max = 172800. ;
  		tilt_time:calendar = "proleptic_gregorian" ;
  		tilt_time:_FillValue = -32767. ;
  		tilt_time:units = "seconds since 2024-07-01" ;
  		tilt_time:valid_min = 0. ;
  	float tilt(tilt_time) ;
  		tilt:_FillValue = -32767.f ;
  		tilt:long_name = "Tilt angle" ;
  		tilt:valid_min = -20.1f ;
  		tilt:valid_max = 20.1f ;
  		tilt:units = "degrees" ;
  	ubyte tilt_flag(tilt_time) ;
  		tilt_flag:_FillValue = 255UB ;
  		tilt_flag:long_name = "Tilt quality flag" ;
  		tilt_flag:flag_values = 0UB, 1UB ;
  		tilt_flag:flag_meanings = "Valid Not_initialized" ;
  	int64 coverage_quality ;
  		coverage_quality:long_name = "coverage quality of navigation data" ;
  		coverage_quality:standard_name = "status_flag" ;
  		coverage_quality:valid_range = 0US, 15US ;
  		coverage_quality:flag_values = 0US, 1US, 2US, 4US, 8US ;
  		coverage_quality:flag_meanings = "good missing-samples too_short_extends no_extend_at_start no_extend_at_end" ;

  // group attributes:
  		:time_coverage_start = "2024-07-01T05:52:23.564Z" ;
  		:time_coverage_end = "2024-07-01T06:48:28.562Z" ;
  } // group navigation_data
}
